library IEEE;
use IEEE.std_logic_1164.all;
--Additional standard or custom libraries go here
package calc_const is
constant DIN1_WIDTH : natural := 16;
constant DIN2_WIDTH : natural := 8;
constant OP_WIDTH : natural := 2;
constant DOUT_WIDTH : natural := 24;
--Other constants, types, subroutines, components go here
end package calc_const;
package body calc_const is
--Subroutine declarations go here
-- you will not have any need for it now, this package is only for defining -
-- some useful constants
end package body calc_const;