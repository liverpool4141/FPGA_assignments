library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use WORK.quantize.all;

package parameters is

--constants
constant pi		:real 		:= 3.14159265359;
constant adc_rate	:integer	:= 64000000;
constant usrp_decim	:integer	:= 250;
constant quad_rate	:integer	:= adc_rate/usrp_decim;
constant audio_decim	:integer	:= 8;
constant audio_rate	:integer	:= quad_rate/audio_decim;
constant volume_level	:integer	:= quantize_f(1.0);
constant samples	:integer	:= 65536*4;
constant audio_samples	:integer 	:= samples/audio_decim;
constant max_taps	:integer	:= 32;
constant max_dev	:real		:= 55000.0;
constant fm_demod_gain	:integer	:= quantize_f(real(quad_rate)/(2.0*pi*max_dev));
constant tau		:real		:= 0.000075;
constant w_pp		:real		:= 0.21140067;

type int_array		is array (integer range <>) of integer;
type char_array	is array (integer range <>) of std_logic_vector(7 downto 0);

--Deemphasis IIR Filter Coefficients:
constant iir_coeff_taps	:integer	:= 2;
constant iir_y_coeffs	:int_array (0 to 1) :=(quantize_f(0.0),quantize_f((w_pp-1.0)/(w_pp+1.0)));
constant iir_x_coeffs	:int_array (0 to 1) :=(quantize_f(w_pp/(1.0+w_pp)),quantize_f(w_pp/(1.0+w_pp)));

--Channel low_pass complex filter coefficients @ 0khz to 80kHz
constant channel_coeff_taps	:integer	:= 20;
constant channel_coeffs_real	:int_array (0 to 19) := (1, 8, -13, 9, 11, -45, 69, -45, -79, 599, 599, -79, -45, 69, -45, 11, 9, -13, 8, 1);
constant channel_coeffs_imag	:int_array (0 to 19)	:= (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0);

--L+R low-pass filter coefficients @15kHz
constant audio_lpr_coeff_taps	:integer	:= 32;
constant audio_lpr_coeffs		:int_array (0 to 31)	:=(-3, -6, -12, -19, -27, -33, -30, -13, 21, 78, 155, 249, 349, 446, 526, 579, 579, 526, 446, 349, 249, 155, 78, 21, -13, -30, -33, -27, -19, -12, -6, -3);

--L-R low-pass filter coefficients @ 15kHz, gain=60
constant audio_lmr_coeff_taps	:integer :=32;
constant audio_lmr_coeffs		:int_array (0 to 31)	:= (-3, -6, -12, -19, -27, -33, -30, -13, 21, 78, 155, 249, 349, 446, 526, 579, 579, 526, 446, 349, 249, 155, 78, 21, -13, -30, -33, -27, -19, -12, -6, -3);

--Pilot tone band-pass filter @ 19kHz
constant bp_pilot_coeff_taps	:integer :=32;
constant bp_pilot_coeffs		:int_array (0 to 31) := (14, 31, 52, 72, 78, 54, -8, -104, -211, -294, -317, -258, -118, 74, 271, 417, 417, 271, 74, -118, -258, -317, -294, -211, -104, -8, 54, 78, 72, 52, 31, 14);

--L-R band-pass filter @ 23kHz to 53kHz
constant bp_lmr_coeff_taps		:integer := 32;
constant bp_lmr_coeffs			:int_array (0 to 31) :=(0, 0, -4, -7, -2, 8, 12, 2, 3, 30, 48, -4, -116, -168, -61, 138, 138, -61, -168, -116, -4, 48, 30, 3, 2, 12, 8, -2, -7, -4, 0, 0);	

--high pass filter @ 0Hz removes noise after pilot tone is squard
constant hp_coeff_taps		:integer	:= 32;
constant hp_coeffs			:int_array (0 to 31) :=(-1, 0, 0, 2, 4, 8, 11, 12, 8, -1, -18, -41, -69, -97, -121, -138, -138, -121, -97, -69, -41, -18, -1, 8, 12, 11, 8, 4, 2, 0, 0, -1);																

constant sin_lut				:int_array (0 to 1023) := (0, 6, 12, 18, 25, 31, 37, 43, 50, 56, 62, 69, 75, 81, 87, 94, 100, 106, 112, 119, 125, 131, 137, 144, 150, 156, 162, 168, 175, 181, 
																187, 193, 199, 205, 212, 218, 224, 230, 236, 242, 248, 254, 260, 267, 273, 279, 285, 291, 297, 303, 309, 315, 321, 327, 333, 339, 344, 350, 
																356, 362, 368, 374, 380, 386, 391, 397, 403, 409, 414, 420, 426, 432, 437, 443, 449, 454, 460, 466, 471, 477, 482, 488, 493, 499, 504, 510, 
																515, 521, 526, 531, 537, 542, 547, 553, 558, 563, 568, 574, 579, 584, 589, 594, 599, 604, 609, 615, 620, 625, 629, 634, 639, 644, 649, 654, 
																659, 664, 668, 673, 678, 683, 687, 692, 696, 701, 706, 710, 715, 719, 724, 728, 732, 737, 741, 745, 750, 754, 758, 762, 767, 771, 775, 779, 
																783, 787, 791, 795, 799, 803, 807, 811, 814, 818, 822, 826, 829, 833, 837, 840, 844, 847, 851, 854, 858, 861, 865, 868, 871, 875, 878, 881, 
																884, 887, 890, 894, 897, 900, 903, 906, 908, 911, 914, 917, 920, 922, 925, 928, 930, 933, 936, 938, 941, 943, 946, 948, 950, 953, 955, 957, 
																959, 962, 964, 966, 968, 970, 972, 974, 976, 978, 979, 981, 983, 985, 986, 988, 990, 991, 993, 994, 996, 997, 999, 1000, 1001, 1003, 1004, 
																1005, 1006, 1007, 1008, 1009, 1010, 1011, 1012, 1013, 1014, 1015, 1016, 1017, 1017, 1018, 1019, 1019, 1020, 1020, 1021, 1021, 1022, 1022, 
																1022, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1023, 1022, 1022, 1022, 1021, 1021, 1020, 1020, 
																1019, 1019, 1018, 1017, 1017, 1016, 1015, 1014, 1013, 1012, 1011, 1010, 1009, 1008, 1007, 1006, 1005, 1004, 1003, 1001, 1000, 999, 997, 996, 
																994, 993, 991, 990, 988, 986, 985, 983, 981, 979, 978, 976, 974, 972, 970, 968, 966, 964, 962, 959, 957, 955, 953, 950, 948, 946, 943, 941, 
																938, 936, 933, 930, 928, 925, 922, 920, 917, 914, 911, 908, 906, 903, 900, 897, 894, 890, 887, 884, 881, 878, 875, 871, 868, 865, 861, 858, 
																854, 851, 847, 844, 840, 837, 833, 829, 826, 822, 818, 814, 811, 807, 803, 799, 795, 791, 787, 783, 779, 775, 771, 767, 762, 758, 754, 750, 
																745, 741, 737, 732, 728, 724, 719, 715, 710, 706, 701, 696, 692, 687, 683, 678, 673, 668, 664, 659, 654, 649, 644, 639, 634, 629, 625, 620, 
																615, 609, 604, 599, 594, 589, 584, 579, 574, 568, 563, 558, 553, 547, 542, 537, 531, 526, 521, 515, 510, 504, 499, 493, 488, 482, 477, 471, 
																466, 460, 454, 449, 443, 437, 432, 426, 420, 414, 409, 403, 397, 391, 386, 380, 374, 368, 362, 356, 350, 344, 339, 333, 327, 321, 315, 309, 
																303, 297, 291, 285, 279, 273, 267, 260, 254, 248, 242, 236, 230, 224, 218, 212, 205, 199, 193, 187, 181, 175, 168, 162, 156, 150, 144, 137, 
																131, 125, 119, 112, 106, 100, 94, 87, 81, 75, 69, 62, 56, 50, 43, 37, 31, 25, 18, 12, 6, 0, -6, -12, -18, -25, -31, -37, -43, -50, -56, -62, 
																-69, -75, -81, -87, -94, -100, -106, -112, -119, -125, -131, -137, -144, -150, -156, -162, -168, -175, -181, -187, -193, -199, -205, -212, 
																-218, -224, -230, -236, -242, -248, -254, -260, -267, -273, -279, -285, -291, -297, -303, -309, -315, -321, -327, -333, -339, -344, -350, 
																-356, -362, -368, -374, -380, -386, -391, -397, -403, -409, -414, -420, -426, -432, -437, -443, -449, -454, -460, -466, -471, -477, -482, 
																-488, -493, -499, -504, -510, -515, -521, -526, -531, -537, -542, -547, -553, -558, -563, -568, -574, -579, -584, -589, -594, -599, -604,
																-609, -615, -620, -625, -629, -634, -639, -644, -649, -654, -659, -664, -668, -673, -678, -683, -687, -692, -696, -701, -706, -710, -715, 
																-719, -724, -728, -732, -737, -741, -745, -750, -754, -758, -762, -767, -771, -775, -779, -783, -787, -791, -795, -799, -803, -807, -811, 
																-814, -818, -822, -826, -829, -833, -837, -840, -844, -847, -851, -854, -858, -861, -865, -868, -871, -875, -878, -881, -884, -887, -890, 
																-894, -897, -900, -903, -906, -908, -911, -914, -917, -920, -922, -925, -928, -930, -933, -936, -938, -941, -943, -946, -948, -950, -953, 
																-955, -957, -959, -962, -964, -966, -968, -970, -972, -974, -976, -978, -979, -981, -983, -985, -986, -988, -990, -991, -993, -994, -996, 
																-997, -999, -1000, -1001, -1003, -1004, -1005, -1006, -1007, -1008, -1009, -1010, -1011, -1012, -1013, -1014, -1015, -1016, -1017, -1017, 
																-1018, -1019, -1019, -1020, -1020, -1021, -1021, -1022, -1022, -1022, -1023, -1023, -1023, -1023, -1023, -1023, -1023, -1023, -1023, -1023, 
																-1023, -1023, -1023, -1023, -1023, -1022, -1022, -1022, -1021, -1021, -1020, -1020, -1019, -1019, -1018, -1017, -1017, -1016, -1015, -1014, 
																-1013, -1012, -1011, -1010, -1009, -1008, -1007, -1006, -1005, -1004, -1003, -1001, -1000, -999, -997, -996, -994, -993, -991, -990, -988, 
																-986, -985, -983, -981, -979, -978, -976, -974, -972, -970, -968, -966, -964, -962, -959, -957, -955, -953, -950, -948, -946, -943, -941, 
																-938, -936, -933, -930, -928, -925, -922, -920, -917, -914, -911, -908, -906, -903, -900, -897, -894, -890, -887, -884, -881, -878, -875, 
																-871, -868, -865, -861, -858, -854, -851, -847, -844, -840, -837, -833, -829, -826, -822, -818, -814, -811, -807, -803, -799, -795, -791,
																-787, -783, -779, -775, -771, -767, -762, -758, -754, -750, -745, -741, -737, -732, -728, -724, -719, -715, -710, -706, -701, -696, -692, 
																-687, -683, -678, -673, -668, -664, -659, -654, -649, -644, -639, -634, -629, -625, -620, -615, -609, -604, -599, -594, -589, -584, -579,
																-574, -568, -563, -558, -553, -547, -542, -537, -531, -526, -521, -515, -510, -504, -499, -493, -488, -482, -477, -471, -466, -460, -454, 
																-449, -443, -437, -432, -426, -420, -414, -409, -403, -397, -391, -386, -380, -374, -368, -362, -356, -350, -344, -339, -333, -327, -321, 
																-315, -309, -303, -297, -291, -285, -279, -273, -267, -260, -254, -248, -242, -236, -230, -224, -218, -212, -205, -199, -193, -187, -181, 
																-175, -168, -162, -156, -150, -144, -137, -131, -125, -119, -112, -106, -100, -94, -87, -81, -75, -69, -62, -56, -50, -43, -37, -31, -25, -18, -12, -6);

end package;



package body parameters is


	
end package body;
